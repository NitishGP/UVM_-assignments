
class apb_sqr extends uvm_sequencer#(apb_tx);
	`uvm_component_utils(apb_sqr)
	`new_component

	
endclass