
class apb_sequencer extends uvm_sequencer#(apb_tx);
  `uvm_component_utils(apb_sequencer)
  `NEW
endclass