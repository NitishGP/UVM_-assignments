
class apb_consumer extends uvm_component;
	`uvm_component_utils(apb_consumer)
	`NEW
	
	function void build_phase(uvm_phase phase);
		super.build_phase(phase);
	endfunction

endclass
