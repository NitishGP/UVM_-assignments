`include "uvm_pkg.sv"
import uvm_pkg::*;

`include "apb_config.sv"
`include "apb_tx.sv"
`include "apb_driver.sv"
`include "apb_stimulus.sv"
`include "apb_convertor.sv"
`include "apb_producer.sv"
`include "apb_consumer.sv"
`include "apb_env.sv"
`include "test_lib.sv"
`include "top.sv"
