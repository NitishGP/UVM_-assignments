
class ahb_base_sequence extends uvm_sequence#(ahb_tx);
	`uvm_object_utils(ahb_base_sequence)
	uvm_phase phase;

	`NEW_OBJ
	
	task pre_body();
		
		uvm_report_info(   "BASE_SQR_SEQ_SEVERITY","INFO FROM BASE SEQ WITH LOW VERBOSITY",UVM_LOW);
		uvm_report_error("BASE_SQR_SEQ_SEVERITY","ERROR FROM BASE SEQ WITH HIGH VERBOSITY",UVM_HIGH);
		uvm_report_warning("BASE_SQR_SEQ_SEVERITY","WARNING FROM BASE SEQ WITH MEDIUM VERBOSITY",UVM_MEDIUM);
		uvm_report_fatal("BASE_SQR_SEQ_SEVERITY","FATAL ERROR MESSAGE FROM Base Seq having verbosity of DEBUG",UVM_DEBUG);


		`uvm_info("BASE_SEQ_PRE_BODY","INSIDE BASE_SEQ_PRE_BODY",UVM_HIGH)
		phase=get_starting_phase();
		if(phase!=null) begin
			phase.raise_objection(null);
		end
	endtask : pre_body

	task body();
		`uvm_info("BASE_SEQ_BODY","INSIDE BASE_SEQ_BODY",UVM_HIGH)
		#10;
		`uvm_do(req);
	endtask : body

	task post_body();
		`uvm_info("BASE_SEQ_POST_BODY","INSIDE BASE_SEQ_POST_BODY",UVM_HIGH)
		if(phase!=null) begin
			phase.drop_objection(null);
		end
	endtask : post_body
endclass : ahb_base_sequence
