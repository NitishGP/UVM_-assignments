module top;
	initial begin
		run_test("apb_base_test");
	end
endmodule
