interface sample_interface(input bit clk,rst);
endinterface
