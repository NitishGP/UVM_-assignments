`include "uvm_macros.svh"
import uvm_pkg::*;

`include "apb_config.sv"
`include "apb_tx.sv"
`include "apb_intf.sv"
`include "apb_seq_lib.sv"
`include "apb_sequencer.sv"
`include "apb_driver.sv"
`include "apb_monitor.sv"
`include "apb_coverage.sv"
`include "apb_agent.sv"
`include "apb_env.sv"
`include "test_lib.sv"
`include "top.sv"