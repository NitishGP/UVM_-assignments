
class sample_tx extends uvm_sequence_item;
	
endclass
