// Code your testbench here
// or browse Examples
`include "list.svh"
