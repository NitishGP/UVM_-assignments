`include "uvm_pkg.sv"
import uvm_pkg::*;


`include "apb_common.sv"
`include "apb_interface.sv"
`include "apb_rtl.v"
`include "apb_tx.sv"
`include "apb_seq_lib.sv"
`include "apb_sqr.sv"
`include "apb_drv.sv"
`include "apb_mon.sv"
`include "apb_cov.sv"
`include "apb_agent.sv"
`include "apb_sbd.sv"
`include "apb_env.sv"
`include "apb_test_lib.sv"
`include "top.sv"
